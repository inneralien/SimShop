/*
    Minimum required tasks for SimShop
*/

// Error reporting
`define report_error         test_util.report_error

// Other conveniences
//`define reset_chip           tb.chip_reset(10)
`define reset_chip           
`define simulation_finish    test_util.simulation_finish
